`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11/18/2020 10:40:29 PM
// Design Name: 
// Module Name: obstacle_rom
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module obstacle_rom(
        input wire clk,
		input wire [4:0] row,
		input wire [4:0] col,
		output reg [11:0] color_data
    );
    (* rom_style = "block" *)

	//signal declaration
	reg [4:0] row_reg;
	reg [4:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @*
	   case ({row_reg, col_reg}) // brick wall skin
	   
	       10'b0000001001: color_data = 12'b111111111111;//9
	       10'b0000010011: color_data = 12'b111111111111;//19
	       
	       10'b0000101001: color_data = 12'b111111111111;//9
	       10'b0000110011: color_data = 12'b111111111111;//19
	       
	       10'b0001001001: color_data = 12'b111111111111;//9
	       10'b0001010011: color_data = 12'b111111111111;//19
	       
	       10'b0001101001: color_data = 12'b111111111111;//9
	       10'b0001110011: color_data = 12'b111111111111;//19
	       
	       10'b0010001001: color_data = 12'b111111111111;//9
	       10'b0010010011: color_data = 12'b111111111111;//19
	       
	       10'b0010100000: color_data = 12'b111111111111;//0
	       10'b0010100001: color_data = 12'b111111111111;//1
	       10'b0010100010: color_data = 12'b111111111111;//2
	       10'b0010100011: color_data = 12'b111111111111;//3
	       10'b0010100100: color_data = 12'b111111111111;//4
	       10'b0010100101: color_data = 12'b111111111111;//5
	       10'b0010100110: color_data = 12'b111111111111;//6
	       10'b0010100111: color_data = 12'b111111111111;//7
	       10'b0010101000: color_data = 12'b111111111111;//8
	       10'b0010101001: color_data = 12'b111111111111;//9
	       10'b0010101010: color_data = 12'b111111111111;//10
	       10'b0010101011: color_data = 12'b111111111111;//11
	       10'b0010101100: color_data = 12'b111111111111;//12
	       10'b0010101101: color_data = 12'b111111111111;//13
	       10'b0010101110: color_data = 12'b111111111111;//14
	       10'b0010101111: color_data = 12'b111111111111;//15
	       10'b0010110000: color_data = 12'b111111111111;//16
	       10'b0010110001: color_data = 12'b111111111111;//17
	       10'b0010110010: color_data = 12'b111111111111;//18
	       10'b0010110011: color_data = 12'b111111111111;//19
	       10'b0010110100: color_data = 12'b111111111111;//20
	       10'b0010110101: color_data = 12'b111111111111;//21
	       10'b0010110110: color_data = 12'b111111111111;//22
	       10'b0010110111: color_data = 12'b111111111111;//23
	       10'b0010111000: color_data = 12'b111111111111;//24
	       10'b0010111001: color_data = 12'b111111111111;//25
	       10'b0010111010: color_data = 12'b111111111111;//26
	       10'b0010111011: color_data = 12'b111111111111;//27
	       10'b0010111100: color_data = 12'b111111111111;//28
	       
	       10'b0011000100: color_data = 12'b111111111111;//4
	       10'b0011001110: color_data = 12'b111111111111;//14
	       10'b0011011000: color_data = 12'b111111111111;//24
	       
	       10'b0011100100: color_data = 12'b111111111111;//4
	       10'b0011101110: color_data = 12'b111111111111;//14
	       10'b0011111000: color_data = 12'b111111111111;//24
	       
	       10'b0100000100: color_data = 12'b111111111111;//4
	       10'b0100001110: color_data = 12'b111111111111;//14
	       10'b0100011000: color_data = 12'b111111111111;//24
	       
	       10'b0100100100: color_data = 12'b111111111111;//4
	       10'b0100101110: color_data = 12'b111111111111;//14
	       10'b0100111000: color_data = 12'b111111111111;//24
	       
	       10'b0101000100: color_data = 12'b111111111111;//4
	       10'b0101001110: color_data = 12'b111111111111;//14
	       10'b0101011000: color_data = 12'b111111111111;//24
	       
	       10'b0101100000: color_data = 12'b111111111111;//0
	       10'b0101100001: color_data = 12'b111111111111;//1
	       10'b0101100010: color_data = 12'b111111111111;//2
	       10'b0101100011: color_data = 12'b111111111111;//3
	       10'b0101100100: color_data = 12'b111111111111;//4
	       10'b0101100101: color_data = 12'b111111111111;//5
	       10'b0101100110: color_data = 12'b111111111111;//6
	       10'b0101100111: color_data = 12'b111111111111;//7
	       10'b0101101000: color_data = 12'b111111111111;//8
	       10'b0101101001: color_data = 12'b111111111111;//9
	       10'b0101101010: color_data = 12'b111111111111;//10
	       10'b0101101011: color_data = 12'b111111111111;//11
	       10'b0101101100: color_data = 12'b111111111111;//12
	       10'b0101101101: color_data = 12'b111111111111;//13
	       10'b0101101110: color_data = 12'b111111111111;//14
	       10'b0101101111: color_data = 12'b111111111111;//15
	       10'b0101110000: color_data = 12'b111111111111;//16
	       10'b0101110001: color_data = 12'b111111111111;//17
	       10'b0101110010: color_data = 12'b111111111111;//18
	       10'b0101110011: color_data = 12'b111111111111;//19
	       10'b0101110100: color_data = 12'b111111111111;//20
	       10'b0101110101: color_data = 12'b111111111111;//21
	       10'b0101110110: color_data = 12'b111111111111;//22
	       10'b0101110111: color_data = 12'b111111111111;//23
	       10'b0101111000: color_data = 12'b111111111111;//24
	       10'b0101111001: color_data = 12'b111111111111;//25
	       10'b0101111010: color_data = 12'b111111111111;//26
	       10'b0101111011: color_data = 12'b111111111111;//27
	       10'b0101111100: color_data = 12'b111111111111;//28
	       
	       10'b0110001001: color_data = 12'b111111111111;//9
	       10'b0110010011: color_data = 12'b111111111111;//19
	       
	       10'b0110101001: color_data = 12'b111111111111;//9
	       10'b0110110011: color_data = 12'b111111111111;//19
	       
	       10'b0111001001: color_data = 12'b111111111111;//9
	       10'b0111010011: color_data = 12'b111111111111;//19
	       
	       10'b0111101001: color_data = 12'b111111111111;//9
	       10'b0111110011: color_data = 12'b111111111111;//19
	       
	       10'b1000001001: color_data = 12'b111111111111;//9
	       10'b1000010011: color_data = 12'b111111111111;//19
	       
	       10'b1000100000: color_data = 12'b111111111111;//0
	       10'b1000100001: color_data = 12'b111111111111;//1
	       10'b1000100010: color_data = 12'b111111111111;//2
	       10'b1000100011: color_data = 12'b111111111111;//3
	       10'b1000100100: color_data = 12'b111111111111;//4
	       10'b1000100101: color_data = 12'b111111111111;//5
	       10'b1000100110: color_data = 12'b111111111111;//6
	       10'b1000100111: color_data = 12'b111111111111;//7
	       10'b1000101000: color_data = 12'b111111111111;//8
	       10'b1000101001: color_data = 12'b111111111111;//9
	       10'b1000101010: color_data = 12'b111111111111;//10
	       10'b1000101011: color_data = 12'b111111111111;//11
	       10'b1000101100: color_data = 12'b111111111111;//12
	       10'b1000101101: color_data = 12'b111111111111;//13
	       10'b1000101110: color_data = 12'b111111111111;//14
	       10'b1000101111: color_data = 12'b111111111111;//15
	       10'b1000110000: color_data = 12'b111111111111;//16
	       10'b1000110001: color_data = 12'b111111111111;//17
	       10'b1000110010: color_data = 12'b111111111111;//18
	       10'b1000110011: color_data = 12'b111111111111;//19
	       10'b1000110100: color_data = 12'b111111111111;//20
	       10'b1000110101: color_data = 12'b111111111111;//21
	       10'b1000110110: color_data = 12'b111111111111;//22
	       10'b1000110111: color_data = 12'b111111111111;//23
	       10'b1000111000: color_data = 12'b111111111111;//24
	       10'b1000111001: color_data = 12'b111111111111;//25
	       10'b1000111010: color_data = 12'b111111111111;//26
	       10'b1000111011: color_data = 12'b111111111111;//27
	       10'b1000111100: color_data = 12'b111111111111;//28
	       
	       10'b1001000100: color_data = 12'b111111111111;//4
	       10'b1001001110: color_data = 12'b111111111111;//14
	       10'b1001011000: color_data = 12'b111111111111;//24
	       
	       10'b1001100100: color_data = 12'b111111111111;//4
	       10'b1001101110: color_data = 12'b111111111111;//14
	       10'b1001111000: color_data = 12'b111111111111;//24
	       
	       10'b1010000100: color_data = 12'b111111111111;//4
	       10'b1010001110: color_data = 12'b111111111111;//14
	       10'b1010011000: color_data = 12'b111111111111;//24
	       
	       10'b1010100100: color_data = 12'b111111111111;//4
	       10'b1010101110: color_data = 12'b111111111111;//14
	       10'b1010111000: color_data = 12'b111111111111;//24
	       
	       10'b1011000100: color_data = 12'b111111111111;//4
	       10'b1011001110: color_data = 12'b111111111111;//14
	       10'b1011011000: color_data = 12'b111111111111;//24
	       
	       10'b1011100000: color_data = 12'b111111111111;//0
	       10'b1011100001: color_data = 12'b111111111111;//1
	       10'b1011100010: color_data = 12'b111111111111;//2
	       10'b1011100011: color_data = 12'b111111111111;//3
	       10'b1011100100: color_data = 12'b111111111111;//4
	       10'b1011100101: color_data = 12'b111111111111;//5
	       10'b1011100110: color_data = 12'b111111111111;//6
	       10'b1011100111: color_data = 12'b111111111111;//7
	       10'b1011101000: color_data = 12'b111111111111;//8
	       10'b1011101001: color_data = 12'b111111111111;//9
	       10'b1011101010: color_data = 12'b111111111111;//10
	       10'b1011101011: color_data = 12'b111111111111;//11
	       10'b1011101100: color_data = 12'b111111111111;//12
	       10'b1011101101: color_data = 12'b111111111111;//13
	       10'b1011101110: color_data = 12'b111111111111;//14
	       10'b1011101111: color_data = 12'b111111111111;//15
	       10'b1011110000: color_data = 12'b111111111111;//16
	       10'b1011110001: color_data = 12'b111111111111;//17
	       10'b1011110010: color_data = 12'b111111111111;//18
	       10'b1011110011: color_data = 12'b111111111111;//19
	       10'b1011110100: color_data = 12'b111111111111;//20
	       10'b1011110101: color_data = 12'b111111111111;//21
	       10'b1011110110: color_data = 12'b111111111111;//22
	       10'b1011110111: color_data = 12'b111111111111;//23
	       10'b1011111000: color_data = 12'b111111111111;//24
	       10'b1011111001: color_data = 12'b111111111111;//25
	       10'b1011111010: color_data = 12'b111111111111;//26
	       10'b1011111011: color_data = 12'b111111111111;//27
	       10'b1011111100: color_data = 12'b111111111111;//28
	       
	       10'b1100001001: color_data = 12'b111111111111;//9
	       10'b1100010011: color_data = 12'b111111111111;//19
	       
	       10'b1100101001: color_data = 12'b111111111111;//9
	       10'b1100110011: color_data = 12'b111111111111;//19
	       
	       10'b1101001001: color_data = 12'b111111111111;//9
	       10'b1101010011: color_data = 12'b111111111111;//19
	       
	       10'b1101101001: color_data = 12'b111111111111;//9
	       10'b1101110011: color_data = 12'b111111111111;//19
	       
	       10'b1110001001: color_data = 12'b111111111111;//9
	       10'b1110010011: color_data = 12'b111111111111;//19
	       
	       10'b1110101001: color_data = 12'b111111111111;//9
	       10'b1110110011: color_data = 12'b111111111111;//19
	       
	       10'b1111000000: color_data = 12'b111111111111;//0
	       10'b1111000001: color_data = 12'b111111111111;//1
	       10'b1111000010: color_data = 12'b111111111111;//2
	       10'b1111000011: color_data = 12'b111111111111;//3
	       10'b1111000100: color_data = 12'b111111111111;//4
	       10'b1111000101: color_data = 12'b111111111111;//5
	       10'b1111000110: color_data = 12'b111111111111;//6
	       10'b1111000111: color_data = 12'b111111111111;//7
	       10'b1111001000: color_data = 12'b111111111111;//8
	       10'b1111001001: color_data = 12'b111111111111;//9
	       10'b1111001010: color_data = 12'b111111111111;//10
	       10'b1111001011: color_data = 12'b111111111111;//11
	       10'b1111001100: color_data = 12'b111111111111;//12
	       10'b1111001101: color_data = 12'b111111111111;//13
	       10'b1111001110: color_data = 12'b111111111111;//14
	       10'b1111001111: color_data = 12'b111111111111;//15
	       10'b1111010000: color_data = 12'b111111111111;//16
	       10'b1111010001: color_data = 12'b111111111111;//17
	       10'b1111010010: color_data = 12'b111111111111;//18
	       10'b1111010011: color_data = 12'b111111111111;//19
	       10'b1111010100: color_data = 12'b111111111111;//20
	       10'b1111010101: color_data = 12'b111111111111;//21
	       10'b1111010110: color_data = 12'b111111111111;//22
	       10'b1111010111: color_data = 12'b111111111111;//23
	       10'b1111011000: color_data = 12'b111111111111;//24
	       10'b1111011001: color_data = 12'b111111111111;//25
	       10'b1111011010: color_data = 12'b111111111111;//26
	       10'b1111011011: color_data = 12'b111111111111;//27
	       10'b1111011100: color_data = 12'b111111111111;//28
	       
	       10'b1111101001: color_data = 12'b111111111111;//9
	       10'b1111110011: color_data = 12'b111111111111;//19
	       
	       default: color_data = 12'b0;
	   endcase
	   
endmodule
