`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11/20/2020 02:37:50 AM
// Design Name: 
// Module Name: space_background
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module space_background(
        input wire clk,
		input wire [8:0] row,
		input wire [9:0] col,
		output reg [11:0] color_data
	);

	(* rom_style = "block" *)

	//signal declaration
	reg [8:0] row_reg;
	reg [9:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @*
	case ({row_reg, col_reg})
	
19'b0001001110011101010: color_data = 12'b111111111111;
19'b0001001110011101011: color_data = 12'b111111111111;
19'b0001010000011101010: color_data = 12'b111111111111;
19'b0001010000011101011: color_data = 12'b111111111111;
19'b0001010010011101010: color_data = 12'b111111111111;
19'b0001010010011101011: color_data = 12'b111111111111;
19'b0001100101000010010: color_data = 12'b111111111111;
19'b0001100101000010011: color_data = 12'b111111111111;
19'b0001100111000010010: color_data = 12'b111111111111;
19'b0001100111000010011: color_data = 12'b111111111111;
19'b0001100111000010100: color_data = 12'b111111111111;
19'b0001101001000010010: color_data = 12'b111111111111;
19'b0001101001000010011: color_data = 12'b111111111111;
19'b0001111000101100101: color_data = 12'b111111111111;
19'b0001111000101100110: color_data = 12'b111111111111;
19'b0001111010001100100: color_data = 12'b111111111111;
19'b0001111010001100101: color_data = 12'b111111111111;
19'b0001111010001100110: color_data = 12'b111111111111;
19'b0001111010001100111: color_data = 12'b111111111111;
19'b0001111010001101000: color_data = 12'b111111111111;
19'b0001111010001101001: color_data = 12'b111111111111;
19'b0001111010101100101: color_data = 12'b111111111111;
19'b0001111010101100110: color_data = 12'b111111111111;
19'b0001111100001100100: color_data = 12'b111111111111;
19'b0001111100001100101: color_data = 12'b111111111111;
19'b0001111100001100110: color_data = 12'b111111111111;
19'b0001111100001100111: color_data = 12'b111111111111;
19'b0001111100001101000: color_data = 12'b111111111111;
19'b0001111100001101001: color_data = 12'b111111111111;
19'b0001111100101100101: color_data = 12'b111111111111;
19'b0001111100101100110: color_data = 12'b111111111111;
19'b0001111110001100100: color_data = 12'b111111111111;
19'b0001111110001100101: color_data = 12'b111111111111;
19'b0001111110001100110: color_data = 12'b111111111111;
19'b0001111110001100111: color_data = 12'b111111111111;
19'b0001111110001101000: color_data = 12'b111111111111;
19'b0001111110001101001: color_data = 12'b111111111111;
19'b0010000000001100100: color_data = 12'b111111111111;
19'b0010000000001100101: color_data = 12'b111111111111;
19'b0010000000001100110: color_data = 12'b111111111111;
19'b0010000000001100111: color_data = 12'b111111111111;
19'b0010000000001101000: color_data = 12'b111111111111;
19'b0010000000001101001: color_data = 12'b111111111111;
19'b0010000010001100100: color_data = 12'b111111111111;
19'b0010000010001100101: color_data = 12'b111111111111;
19'b0010000010001100110: color_data = 12'b111111111111;
19'b0010000010001100111: color_data = 12'b111111111111;
19'b0010000010001101000: color_data = 12'b111111111111;
19'b0010000010001101001: color_data = 12'b111111111111;
19'b0010000100001100100: color_data = 12'b111111111111;
19'b0010000100001100101: color_data = 12'b111111111111;
19'b0010000100001100110: color_data = 12'b111111111111;
19'b0010000100001100111: color_data = 12'b111111111111;
19'b0010000100001101000: color_data = 12'b111111111111;
19'b0010000100001101001: color_data = 12'b111111111111;
19'b0010011010110110010: color_data = 12'b111111111111;
19'b0010011100110110001: color_data = 12'b111111111111;
19'b0010011100110110010: color_data = 12'b111111111111;
19'b0010011100110110011: color_data = 12'b111111111111;
19'b0010011110110110010: color_data = 12'b111111111111;
19'b0010101111000001001: color_data = 12'b111111111111;
19'b0010110001000001000: color_data = 12'b111111111111;
19'b0010110001000001001: color_data = 12'b111111111111;
19'b0010110001000001010: color_data = 12'b111111111111;
19'b0010110011000001000: color_data = 12'b111111111111;
19'b0010110011000001001: color_data = 12'b111111111111;
19'b0010110011000001010: color_data = 12'b111111111111;
19'b0010111001000111011: color_data = 12'b111111111111;
19'b0010111001000111100: color_data = 12'b111111111111;
19'b0010111001000111101: color_data = 12'b111111111111;
19'b0010111001000111110: color_data = 12'b111111111111;
19'b0010111001000111111: color_data = 12'b111111111111;
19'b0010111001001000000: color_data = 12'b111111111111;
19'b0010111001001000001: color_data = 12'b111111111111;
19'b0010111001001000010: color_data = 12'b111111111111;
19'b0010111001001000011: color_data = 12'b111111111111;
19'b0010111001001000100: color_data = 12'b111111111111;
19'b0010111001001000101: color_data = 12'b111111111111;
19'b0010111001001000110: color_data = 12'b111111111111;
19'b0010111011000111011: color_data = 12'b111111111111;
19'b0010111011000111100: color_data = 12'b111111111111;
19'b0010111011000111101: color_data = 12'b111111111111;
19'b0010111011000111110: color_data = 12'b111111111111;
19'b0010111011000111111: color_data = 12'b111111111111;
19'b0010111011001000000: color_data = 12'b111111111111;
19'b0010111011001000001: color_data = 12'b111111111111;
19'b0010111011001000010: color_data = 12'b111111111111;
19'b0010111011001000011: color_data = 12'b111111111111;
19'b0010111011001000100: color_data = 12'b111111111111;
19'b0010111011001000101: color_data = 12'b111111111111;
19'b0010111011001000110: color_data = 12'b111111111111;
19'b0010111101000111011: color_data = 12'b111111111111;
19'b0010111101000111100: color_data = 12'b111111111111;
19'b0010111101000111101: color_data = 12'b111111111111;
19'b0010111101000111110: color_data = 12'b111111111111;
19'b0010111101000111111: color_data = 12'b111111111111;
19'b0010111101001000000: color_data = 12'b111111111111;
19'b0010111101001000001: color_data = 12'b111111111111;
19'b0010111101001000010: color_data = 12'b111111111111;
19'b0010111101001000011: color_data = 12'b111111111111;
19'b0010111101001000100: color_data = 12'b111111111111;
19'b0010111101001000101: color_data = 12'b111111111111;
19'b0010111101001000110: color_data = 12'b111111111111;
19'b0010111110011001010: color_data = 12'b111111111111;
19'b0010111110011001011: color_data = 12'b111111111111;
19'b0010111111000111011: color_data = 12'b111111111111;
19'b0010111111000111100: color_data = 12'b111111111111;
19'b0010111111000111101: color_data = 12'b111111111111;
19'b0010111111000111110: color_data = 12'b111111111111;
19'b0010111111000111111: color_data = 12'b111111111111;
19'b0010111111001000000: color_data = 12'b111111111111;
19'b0010111111001000001: color_data = 12'b111111111111;
19'b0010111111001000010: color_data = 12'b111111111111;
19'b0010111111001000011: color_data = 12'b111111111111;
19'b0010111111001000100: color_data = 12'b111111111111;
19'b0010111111001000101: color_data = 12'b111111111111;
19'b0010111111001000110: color_data = 12'b111111111111;
19'b0011000000011001010: color_data = 12'b111111111111;
19'b0011000000011001011: color_data = 12'b111111111111;
19'b0011000001000111011: color_data = 12'b111111111111;
19'b0011000001000111100: color_data = 12'b111111111111;
19'b0011000001000111101: color_data = 12'b111111111111;
19'b0011000001000111110: color_data = 12'b111111111111;
19'b0011000001000111111: color_data = 12'b111111111111;
19'b0011000001001000000: color_data = 12'b111111111111;
19'b0011000001001000001: color_data = 12'b111111111111;
19'b0011000001001000010: color_data = 12'b111111111111;
19'b0011000001001000011: color_data = 12'b111111111111;
19'b0011000001001000100: color_data = 12'b111111111111;
19'b0011000001001000101: color_data = 12'b111111111111;
19'b0011000001001000110: color_data = 12'b111111111111;
19'b0011000011000111011: color_data = 12'b111111111111;
19'b0011000011000111100: color_data = 12'b111111111111;
19'b0011000011000111101: color_data = 12'b111111111111;
19'b0011000011000111110: color_data = 12'b111111111111;
19'b0011000011000111111: color_data = 12'b111111111111;
19'b0011000011001000000: color_data = 12'b111111111111;
19'b0011000011001000001: color_data = 12'b111111111111;
19'b0011000011001000010: color_data = 12'b111111111111;
19'b0011000011001000011: color_data = 12'b111111111111;
19'b0011000011001000100: color_data = 12'b111111111111;
19'b0011000011001000101: color_data = 12'b111111111111;
19'b0011000011001000110: color_data = 12'b111111111111;
19'b0011000101000111011: color_data = 12'b111111111111;
19'b0011000101000111100: color_data = 12'b111111111111;
19'b0011000101000111101: color_data = 12'b111111111111;
19'b0011000101000111110: color_data = 12'b111111111111;
19'b0011000101000111111: color_data = 12'b111111111111;
19'b0011000101001000000: color_data = 12'b111111111111;
19'b0011000101001000001: color_data = 12'b111111111111;
19'b0011000101001000010: color_data = 12'b111111111111;
19'b0011000101001000011: color_data = 12'b111111111111;
19'b0011000101001000100: color_data = 12'b111111111111;
19'b0011000101001000101: color_data = 12'b111111111111;
19'b0011000101001000110: color_data = 12'b111111111111;
19'b0011000111000111011: color_data = 12'b111111111111;
19'b0011000111000111100: color_data = 12'b111111111111;
19'b0011000111000111101: color_data = 12'b111111111111;
19'b0011000111000111110: color_data = 12'b111111111111;
19'b0011000111000111111: color_data = 12'b111111111111;
19'b0011000111001000000: color_data = 12'b111111111111;
19'b0011000111001000001: color_data = 12'b111111111111;
19'b0011000111001000010: color_data = 12'b111111111111;
19'b0011000111001000011: color_data = 12'b111111111111;
19'b0011000111001000100: color_data = 12'b111111111111;
19'b0011000111001000101: color_data = 12'b111111111111;
19'b0011000111001000110: color_data = 12'b111111111111;
19'b0011001001000111011: color_data = 12'b111111111111;
19'b0011001001000111100: color_data = 12'b111111111111;
19'b0011001001000111101: color_data = 12'b111111111111;
19'b0011001001000111110: color_data = 12'b111111111111;
19'b0011001001000111111: color_data = 12'b111111111111;
19'b0011001001001000000: color_data = 12'b111111111111;
19'b0011001001001000001: color_data = 12'b111111111111;
19'b0011001001001000010: color_data = 12'b111111111111;
19'b0011001001001000011: color_data = 12'b111111111111;
19'b0011001001001000100: color_data = 12'b111111111111;
19'b0011001001001000101: color_data = 12'b111111111111;
19'b0011001001001000110: color_data = 12'b111111111111;
19'b0011001011000111011: color_data = 12'b111111111111;
19'b0011001011000111100: color_data = 12'b111111111111;
19'b0011001011000111101: color_data = 12'b111111111111;
19'b0011001011000111110: color_data = 12'b111111111111;
19'b0011001011000111111: color_data = 12'b111111111111;
19'b0011001011001000000: color_data = 12'b111111111111;
19'b0011001011001000001: color_data = 12'b111111111111;
19'b0011001011001000010: color_data = 12'b111111111111;
19'b0011001011001000011: color_data = 12'b111111111111;
19'b0011001011001000100: color_data = 12'b111111111111;
19'b0011001011001000101: color_data = 12'b111111111111;
19'b0011001011001000110: color_data = 12'b111111111111;
19'b0011001101000111011: color_data = 12'b111111111111;
19'b0011001101000111100: color_data = 12'b111111111111;
19'b0011001101000111101: color_data = 12'b111111111111;
19'b0011001101000111110: color_data = 12'b111111111111;
19'b0011001101000111111: color_data = 12'b111111111111;
19'b0011001101001000000: color_data = 12'b111111111111;
19'b0011001101001000001: color_data = 12'b111111111111;
19'b0011001101001000010: color_data = 12'b111111111111;
19'b0011001101001000011: color_data = 12'b111111111111;
19'b0011001101001000100: color_data = 12'b111111111111;
19'b0011001101001000101: color_data = 12'b111111111111;
19'b0011001101001000110: color_data = 12'b111111111111;
19'b0011001111000111100: color_data = 12'b111111111111;
19'b0011001111000111101: color_data = 12'b111111111111;
19'b0011001111000111110: color_data = 12'b111111111111;
19'b0011001111000111111: color_data = 12'b111111111111;
19'b0011001111001000000: color_data = 12'b111111111111;
19'b0011001111001000001: color_data = 12'b111111111111;
19'b0011001111001000010: color_data = 12'b111111111111;
19'b0011001111001000011: color_data = 12'b111111111111;
19'b0011001111001000100: color_data = 12'b111111111111;
19'b0011001111001000101: color_data = 12'b111111111111;
19'b0011001111001000110: color_data = 12'b111111111111;
19'b0011111010100011111: color_data = 12'b111111111111;
19'b0011111010100100000: color_data = 12'b111111111111;
19'b0011111100100011111: color_data = 12'b111111111111;
19'b0011111100100100000: color_data = 12'b111111111111;
19'b0100010110010000001: color_data = 12'b111111111111;
19'b0100010110010000010: color_data = 12'b111111111111;
19'b0100010110010000011: color_data = 12'b111111111111;
19'b0100010110010000100: color_data = 12'b111111111111;
19'b0100010110010000101: color_data = 12'b111111111111;
19'b0100010110110010101: color_data = 12'b111111111111;
19'b0100010110110010110: color_data = 12'b111111111111;
19'b0100011000010000001: color_data = 12'b111111111111;
19'b0100011000010000010: color_data = 12'b111111111111;
19'b0100011000010000011: color_data = 12'b111111111111;
19'b0100011000010000100: color_data = 12'b111111111111;
19'b0100011000010000101: color_data = 12'b111111111111;
19'b0100011000110010101: color_data = 12'b111111111111;
19'b0100011000110010110: color_data = 12'b111111111111;
19'b0100011010010000001: color_data = 12'b111111111111;
19'b0100011010010000010: color_data = 12'b111111111111;
19'b0100011010010000011: color_data = 12'b111111111111;
19'b0100011010010000100: color_data = 12'b111111111111;
19'b0100011010010000101: color_data = 12'b111111111111;
19'b0100011100010000001: color_data = 12'b111111111111;
19'b0100011100010000010: color_data = 12'b111111111111;
19'b0100011100010000011: color_data = 12'b111111111111;
19'b0100011100010000100: color_data = 12'b111111111111;
19'b0100011100010000101: color_data = 12'b111111111111;
19'b0100011110010000001: color_data = 12'b111111111111;
19'b0100011110010000010: color_data = 12'b111111111111;
19'b0100011110010000011: color_data = 12'b111111111111;
19'b0100011110010000100: color_data = 12'b111111111111;
19'b0100011110010000101: color_data = 12'b111111111111;
19'b0100110000100011011: color_data = 12'b111111111111;
19'b0100110000100011100: color_data = 12'b111111111111;
19'b0100110010100011011: color_data = 12'b111111111111;
19'b0100110010100011100: color_data = 12'b111111111111;
19'b0100110100111110000: color_data = 12'b111111111111;
19'b0100110100111110001: color_data = 12'b111111111111;
19'b0100110110111110000: color_data = 12'b111111111111;
19'b0100110110111110001: color_data = 12'b111111111111;
19'b0100111000111110000: color_data = 12'b111111111111;
19'b0110000000101011101: color_data = 12'b111111111111;
19'b0110000000101011110: color_data = 12'b111111111111;
19'b0110000000101011111: color_data = 12'b111111111111;
19'b0110000010101011101: color_data = 12'b111111111111;
19'b0110000010101011110: color_data = 12'b111111111111;
19'b0110000010101011111: color_data = 12'b111111111111;
19'b0110000100101011101: color_data = 12'b111111111111;
19'b0110000100101011110: color_data = 12'b111111111111;
19'b0110001100001010011: color_data = 12'b111111111111;
19'b0110001100001010100: color_data = 12'b111111111111;
19'b0110001100001010101: color_data = 12'b111111111111;
19'b0110001110001010011: color_data = 12'b111111111111;
19'b0110001110001010100: color_data = 12'b111111111111;
19'b0110001110001010101: color_data = 12'b111111111111;
19'b0110100000011001001: color_data = 12'b111111111111;
19'b0110100000011001010: color_data = 12'b111111111111;
19'b0110100010011001001: color_data = 12'b111111111111;
19'b0110100010011001010: color_data = 12'b111111111111;
19'b0110100100011001001: color_data = 12'b111111111111;
19'b0110100100011001010: color_data = 12'b111111111111;
19'b0110101010110010001: color_data = 12'b111111111111;
19'b0110101010110010010: color_data = 12'b111111111111;
19'b0110101010110010011: color_data = 12'b111111111111;
19'b0110101010110010100: color_data = 12'b111111111111;
19'b0110101010110010101: color_data = 12'b111111111111;
19'b0110101010110010110: color_data = 12'b111111111111;
19'b0110101100110010001: color_data = 12'b111111111111;
19'b0110101100110010010: color_data = 12'b111111111111;
19'b0110101100110010011: color_data = 12'b111111111111;
19'b0110101100110010100: color_data = 12'b111111111111;
19'b0110101100110010101: color_data = 12'b111111111111;
19'b0110101100110010110: color_data = 12'b111111111111;
19'b0110101110110010001: color_data = 12'b111111111111;
19'b0110101110110010010: color_data = 12'b111111111111;
19'b0110101110110010011: color_data = 12'b111111111111;
19'b0110101110110010100: color_data = 12'b111111111111;
19'b0110101110110010101: color_data = 12'b111111111111;
19'b0110101110110010110: color_data = 12'b111111111111;
19'b0110110000110010001: color_data = 12'b111111111111;
19'b0110110000110010010: color_data = 12'b111111111111;
19'b0110110000110010011: color_data = 12'b111111111111;
19'b0110110000110010100: color_data = 12'b111111111111;
19'b0110110000110010101: color_data = 12'b111111111111;
19'b0110110000110010110: color_data = 12'b111111111111;
19'b0110110010110010001: color_data = 12'b111111111111;
19'b0110110010110010010: color_data = 12'b111111111111;
19'b0110110010110010011: color_data = 12'b111111111111;
19'b0110110010110010100: color_data = 12'b111111111111;
19'b0110110010110010101: color_data = 12'b111111111111;
19'b0110110010110010110: color_data = 12'b111111111111;
19'b0110110100110010001: color_data = 12'b111111111111;
19'b0110110100110010010: color_data = 12'b111111111111;
19'b0110110100110010011: color_data = 12'b111111111111;
19'b0110110100110010100: color_data = 12'b111111111111;
19'b0110110100110010101: color_data = 12'b111111111111;
19'b0110110100110010110: color_data = 12'b111111111111;
19'b0110110110110010001: color_data = 12'b111111111111;
19'b0110110110110010010: color_data = 12'b111111111111;
19'b0110110110110010011: color_data = 12'b111111111111;
19'b0110110110110010100: color_data = 12'b111111111111;
19'b0110110110110010101: color_data = 12'b111111111111;
19'b0110110110110010110: color_data = 12'b111111111111;
19'b0110111001000001011: color_data = 12'b111111111111;
19'b0110111001000001100: color_data = 12'b111111111111;
19'b0110111001000001101: color_data = 12'b111111111111;
19'b0110111010100110010: color_data = 12'b111111111111;
19'b0110111010100110011: color_data = 12'b111111111111;
19'b0110111011000001011: color_data = 12'b111111111111;
19'b0110111011000001100: color_data = 12'b111111111111;
19'b0110111100100110010: color_data = 12'b111111111111;
19'b0110111100100110011: color_data = 12'b111111111111;
19'b0111000100101111001: color_data = 12'b111111111111;
19'b0111000100101111010: color_data = 12'b111111111111;
19'b0111000110101111001: color_data = 12'b111111111111;
19'b0111000110101111010: color_data = 12'b111111111111;
19'b1000100110011111111: color_data = 12'b111111111111;
19'b1000100110100000000: color_data = 12'b111111111111;
19'b1000101000011111110: color_data = 12'b111111111111;
19'b1000101000011111111: color_data = 12'b111111111111;
19'b1000101000100000000: color_data = 12'b111111111111;
19'b1000101001001000101: color_data = 12'b111111111111;
19'b1000101010011111111: color_data = 12'b111111111111;
19'b1000101010100000000: color_data = 12'b111111111111;
19'b1000101011001000100: color_data = 12'b111111111111;
19'b1000101011001000101: color_data = 12'b111111111111;
19'b1000101011001000110: color_data = 12'b111111111111;
19'b1000101101001000100: color_data = 12'b111111111111;
19'b1000101101001000101: color_data = 12'b111111111111;
19'b1000101101001000110: color_data = 12'b111111111111;
19'b1001011110110101111: color_data = 12'b111111111111;
19'b1001011110110110000: color_data = 12'b111111111111;
19'b1001100000110101110: color_data = 12'b111111111111;
19'b1001100000110101111: color_data = 12'b111111111111;
19'b1001100000110110000: color_data = 12'b111111111111;
19'b1001101010000111111: color_data = 12'b111111111111;
19'b1001101010001000000: color_data = 12'b111111111111;
19'b1001101100000111110: color_data = 12'b111111111111;
19'b1001101100000111111: color_data = 12'b111111111111;
19'b1001101100001000000: color_data = 12'b111111111111;
19'b1001101110000111111: color_data = 12'b111111111111;
19'b1001101110001000000: color_data = 12'b111111111111;
19'b1001110000101001100: color_data = 12'b111111111111;
19'b1001110000101001101: color_data = 12'b111111111111;
19'b1001110010101001100: color_data = 12'b111111111111;
19'b1001110010101001101: color_data = 12'b111111111111;
19'b1001110011000111011: color_data = 12'b111111111111;
19'b1001110011000111100: color_data = 12'b111111111111;
19'b1001110101000111011: color_data = 12'b111111111111;
19'b1001110101000111100: color_data = 12'b111111111111;
19'b1001110101000111101: color_data = 12'b111111111111;
19'b1001110111000111011: color_data = 12'b111111111111;
19'b1001110111000111100: color_data = 12'b111111111111;
19'b1001111010001011001: color_data = 12'b111111111111;
19'b1001111010001011010: color_data = 12'b111111111111;
19'b1001111100001011001: color_data = 12'b111111111111;
19'b1001111100001011010: color_data = 12'b111111111111;
19'b1001111110001011001: color_data = 12'b111111111111;
19'b1010010100010011100: color_data = 12'b111111111111;
19'b1010010100010011101: color_data = 12'b111111111111;
19'b1010010100010011110: color_data = 12'b111111111111;
19'b1010010100010011111: color_data = 12'b111111111111;
19'b1010010100010100000: color_data = 12'b111111111111;
19'b1010010100010100001: color_data = 12'b111111111111;
19'b1010010110010011100: color_data = 12'b111111111111;
19'b1010010110010011101: color_data = 12'b111111111111;
19'b1010010110010011110: color_data = 12'b111111111111;
19'b1010010110010011111: color_data = 12'b111111111111;
19'b1010010110010100000: color_data = 12'b111111111111;
19'b1010010110010100001: color_data = 12'b111111111111;
19'b1010011000010011100: color_data = 12'b111111111111;
19'b1010011000010011101: color_data = 12'b111111111111;
19'b1010011000010011110: color_data = 12'b111111111111;
19'b1010011000010011111: color_data = 12'b111111111111;
19'b1010011000010100000: color_data = 12'b111111111111;
19'b1010011000010100001: color_data = 12'b111111111111;
19'b1010011010010011100: color_data = 12'b111111111111;
19'b1010011010010011101: color_data = 12'b111111111111;
19'b1010011010010011110: color_data = 12'b111111111111;
19'b1010011010010011111: color_data = 12'b111111111111;
19'b1010011010010100000: color_data = 12'b111111111111;
19'b1010011010010100001: color_data = 12'b111111111111;
19'b1010011100010011100: color_data = 12'b111111111111;
19'b1010011100010011101: color_data = 12'b111111111111;
19'b1010011100010011110: color_data = 12'b111111111111;
19'b1010011100010011111: color_data = 12'b111111111111;
19'b1010011100010100000: color_data = 12'b111111111111;
19'b1010011100010100001: color_data = 12'b111111111111;
19'b1010011110010011100: color_data = 12'b111111111111;
19'b1010011110010011101: color_data = 12'b111111111111;
19'b1010011110010011110: color_data = 12'b111111111111;
19'b1010011110010011111: color_data = 12'b111111111111;
19'b1010011110010100000: color_data = 12'b111111111111;
19'b1010011110010100001: color_data = 12'b111111111111;
19'b1011101000011111100: color_data = 12'b111111111111;
19'b1011101000011111101: color_data = 12'b111111111111;
19'b1011101010011111100: color_data = 12'b111111111111;
19'b1011101010011111101: color_data = 12'b111111111111;
19'b1011101100011111100: color_data = 12'b111111111111;
19'b1011101100011111101: color_data = 12'b111111111111;
19'b1100000110010001111: color_data = 12'b111111111111;
19'b1100000110010010000: color_data = 12'b111111111111;
19'b1100000110010010001: color_data = 12'b111111111111;
19'b1100001000010010000: color_data = 12'b111111111111;
19'b1100001000010010001: color_data = 12'b111111111111;
19'b1100001000101011000: color_data = 12'b111111111111;
19'b1100001010010010000: color_data = 12'b111111111111;
19'b1100001010010010001: color_data = 12'b111111111111;
19'b1100001010101010111: color_data = 12'b111111111111;
19'b1100001010101011000: color_data = 12'b111111111111;
19'b1100001010101011001: color_data = 12'b111111111111;
19'b1100001011000101110: color_data = 12'b111111111111;
19'b1100001011000101111: color_data = 12'b111111111111;
19'b1100001011000110000: color_data = 12'b111111111111;
19'b1100001100010010000: color_data = 12'b111111111111;
19'b1100001100101011000: color_data = 12'b111111111111;
19'b1100001101000101110: color_data = 12'b111111111111;
19'b1100001101000101111: color_data = 12'b111111111111;
19'b1100001101000110000: color_data = 12'b111111111111;
19'b1100001111000101110: color_data = 12'b111111111111;
19'b1100001111000101111: color_data = 12'b111111111111;
19'b1100001111000110000: color_data = 12'b111111111111;
19'b1100110100110100100: color_data = 12'b111111111111;
19'b1100110100110100101: color_data = 12'b111111111111;
19'b1100110100110100110: color_data = 12'b111111111111;
19'b1100110100110100111: color_data = 12'b111111111111;
19'b1100110100110101000: color_data = 12'b111111111111;
19'b1100110100110101001: color_data = 12'b111111111111;
19'b1100110100110101010: color_data = 12'b111111111111;
19'b1100110100110101011: color_data = 12'b111111111111;
19'b1100110100110101100: color_data = 12'b111111111111;
19'b1100110100110101101: color_data = 12'b111111111111;
19'b1100110100110101110: color_data = 12'b111111111111;
19'b1100110110110100011: color_data = 12'b111111111111;
19'b1100110110110100100: color_data = 12'b111111111111;
19'b1100110110110100101: color_data = 12'b111111111111;
19'b1100110110110100110: color_data = 12'b111111111111;
19'b1100110110110100111: color_data = 12'b111111111111;
19'b1100110110110101000: color_data = 12'b111111111111;
19'b1100110110110101001: color_data = 12'b111111111111;
19'b1100110110110101010: color_data = 12'b111111111111;
19'b1100110110110101011: color_data = 12'b111111111111;
19'b1100110110110101100: color_data = 12'b111111111111;
19'b1100110110110101101: color_data = 12'b111111111111;
19'b1100110110110101110: color_data = 12'b111111111111;
19'b1100111000110100011: color_data = 12'b111111111111;
19'b1100111000110100100: color_data = 12'b111111111111;
19'b1100111000110100101: color_data = 12'b111111111111;
19'b1100111000110100110: color_data = 12'b111111111111;
19'b1100111000110100111: color_data = 12'b111111111111;
19'b1100111000110101000: color_data = 12'b111111111111;
19'b1100111000110101001: color_data = 12'b111111111111;
19'b1100111000110101010: color_data = 12'b111111111111;
19'b1100111000110101011: color_data = 12'b111111111111;
19'b1100111000110101100: color_data = 12'b111111111111;
19'b1100111000110101101: color_data = 12'b111111111111;
19'b1100111000110101110: color_data = 12'b111111111111;
19'b1100111010110100011: color_data = 12'b111111111111;
19'b1100111010110100100: color_data = 12'b111111111111;
19'b1100111010110100101: color_data = 12'b111111111111;
19'b1100111010110100110: color_data = 12'b111111111111;
19'b1100111010110100111: color_data = 12'b111111111111;
19'b1100111010110101000: color_data = 12'b111111111111;
19'b1100111010110101001: color_data = 12'b111111111111;
19'b1100111010110101010: color_data = 12'b111111111111;
19'b1100111010110101011: color_data = 12'b111111111111;
19'b1100111010110101100: color_data = 12'b111111111111;
19'b1100111010110101101: color_data = 12'b111111111111;
19'b1100111010110101110: color_data = 12'b111111111111;
19'b1100111010111111010: color_data = 12'b111111111111;
19'b1100111010111111011: color_data = 12'b111111111111;
19'b1100111100110100011: color_data = 12'b111111111111;
19'b1100111100110100100: color_data = 12'b111111111111;
19'b1100111100110100101: color_data = 12'b111111111111;
19'b1100111100110100110: color_data = 12'b111111111111;
19'b1100111100110100111: color_data = 12'b111111111111;
19'b1100111100110101000: color_data = 12'b111111111111;
19'b1100111100110101001: color_data = 12'b111111111111;
19'b1100111100110101010: color_data = 12'b111111111111;
19'b1100111100110101011: color_data = 12'b111111111111;
19'b1100111100110101100: color_data = 12'b111111111111;
19'b1100111100110101101: color_data = 12'b111111111111;
19'b1100111100110101110: color_data = 12'b111111111111;
19'b1100111100111111010: color_data = 12'b111111111111;
19'b1100111100111111011: color_data = 12'b111111111111;
19'b1100111110110100011: color_data = 12'b111111111111;
19'b1100111110110100100: color_data = 12'b111111111111;
19'b1100111110110100101: color_data = 12'b111111111111;
19'b1100111110110100110: color_data = 12'b111111111111;
19'b1100111110110100111: color_data = 12'b111111111111;
19'b1100111110110101000: color_data = 12'b111111111111;
19'b1100111110110101001: color_data = 12'b111111111111;
19'b1100111110110101010: color_data = 12'b111111111111;
19'b1100111110110101011: color_data = 12'b111111111111;
19'b1100111110110101100: color_data = 12'b111111111111;
19'b1100111110110101101: color_data = 12'b111111111111;
19'b1100111110110101110: color_data = 12'b111111111111;
19'b1100111110111111001: color_data = 12'b111111111111;
19'b1101000000110100011: color_data = 12'b111111111111;
19'b1101000000110100100: color_data = 12'b111111111111;
19'b1101000000110100101: color_data = 12'b111111111111;
19'b1101000000110100110: color_data = 12'b111111111111;
19'b1101000000110100111: color_data = 12'b111111111111;
19'b1101000000110101000: color_data = 12'b111111111111;
19'b1101000000110101001: color_data = 12'b111111111111;
19'b1101000000110101010: color_data = 12'b111111111111;
19'b1101000000110101011: color_data = 12'b111111111111;
19'b1101000000110101100: color_data = 12'b111111111111;
19'b1101000000110101101: color_data = 12'b111111111111;
19'b1101000000110101110: color_data = 12'b111111111111;
19'b1101000010110100011: color_data = 12'b111111111111;
19'b1101000010110100100: color_data = 12'b111111111111;
19'b1101000010110100101: color_data = 12'b111111111111;
19'b1101000010110100110: color_data = 12'b111111111111;
19'b1101000010110100111: color_data = 12'b111111111111;
19'b1101000010110101000: color_data = 12'b111111111111;
19'b1101000010110101001: color_data = 12'b111111111111;
19'b1101000010110101010: color_data = 12'b111111111111;
19'b1101000010110101011: color_data = 12'b111111111111;
19'b1101000010110101100: color_data = 12'b111111111111;
19'b1101000010110101101: color_data = 12'b111111111111;
19'b1101000010110101110: color_data = 12'b111111111111;
19'b1101000100110100011: color_data = 12'b111111111111;
19'b1101000100110100100: color_data = 12'b111111111111;
19'b1101000100110100101: color_data = 12'b111111111111;
19'b1101000100110100110: color_data = 12'b111111111111;
19'b1101000100110100111: color_data = 12'b111111111111;
19'b1101000100110101000: color_data = 12'b111111111111;
19'b1101000100110101001: color_data = 12'b111111111111;
19'b1101000100110101010: color_data = 12'b111111111111;
19'b1101000100110101011: color_data = 12'b111111111111;
19'b1101000100110101100: color_data = 12'b111111111111;
19'b1101000100110101101: color_data = 12'b111111111111;
19'b1101000100110101110: color_data = 12'b111111111111;
19'b1101000110110100011: color_data = 12'b111111111111;
19'b1101000110110100100: color_data = 12'b111111111111;
19'b1101000110110100101: color_data = 12'b111111111111;
19'b1101000110110100110: color_data = 12'b111111111111;
19'b1101000110110100111: color_data = 12'b111111111111;
19'b1101000110110101000: color_data = 12'b111111111111;
19'b1101000110110101001: color_data = 12'b111111111111;
19'b1101000110110101010: color_data = 12'b111111111111;
19'b1101000110110101011: color_data = 12'b111111111111;
19'b1101000110110101100: color_data = 12'b111111111111;
19'b1101000110110101101: color_data = 12'b111111111111;
19'b1101000110110101110: color_data = 12'b111111111111;
19'b1101001000110100011: color_data = 12'b111111111111;
19'b1101001000110100100: color_data = 12'b111111111111;
19'b1101001000110100101: color_data = 12'b111111111111;
19'b1101001000110100110: color_data = 12'b111111111111;
19'b1101001000110100111: color_data = 12'b111111111111;
19'b1101001000110101000: color_data = 12'b111111111111;
19'b1101001000110101001: color_data = 12'b111111111111;
19'b1101001000110101010: color_data = 12'b111111111111;
19'b1101001000110101011: color_data = 12'b111111111111;
19'b1101001000110101100: color_data = 12'b111111111111;
19'b1101001000110101101: color_data = 12'b111111111111;
19'b1101001000110101110: color_data = 12'b111111111111;
19'b1101001010110100011: color_data = 12'b111111111111;
19'b1101001010110100100: color_data = 12'b111111111111;
19'b1101001010110100101: color_data = 12'b111111111111;
19'b1101001010110100110: color_data = 12'b111111111111;
19'b1101001010110100111: color_data = 12'b111111111111;
19'b1101001010110101000: color_data = 12'b111111111111;
19'b1101001010110101001: color_data = 12'b111111111111;
19'b1101001010110101010: color_data = 12'b111111111111;
19'b1101001010110101011: color_data = 12'b111111111111;
19'b1101001010110101100: color_data = 12'b111111111111;
19'b1101001010110101101: color_data = 12'b111111111111;
19'b1101001010110101110: color_data = 12'b111111111111;
19'b1101001100000111010: color_data = 12'b111111111111;
19'b1101001100000111011: color_data = 12'b111111111111;
19'b1101001110000111010: color_data = 12'b111111111111;
19'b1101001110000111011: color_data = 12'b111111111111;
19'b1101100110100001010: color_data = 12'b111111111111;
19'b1101100110100001011: color_data = 12'b111111111111;
19'b1101100110100001100: color_data = 12'b111111111111;
19'b1101101000100001010: color_data = 12'b111111111111;
19'b1101101000100001011: color_data = 12'b111111111111;
19'b1101101000100001100: color_data = 12'b111111111111;
19'b1101101100010101010: color_data = 12'b111111111111;
19'b1101101100010101011: color_data = 12'b111111111111;
19'b1101101110010101010: color_data = 12'b111111111111;
19'b1101101110010101011: color_data = 12'b111111111111;
19'b1101101110010101100: color_data = 12'b111111111111;
19'b1101110000010101010: color_data = 12'b111111111111;
19'b1101110000010101011: color_data = 12'b111111111111;


	   
	   default: color_data = 12'b0;
	endcase
endmodule
